/*
实现彩虹效果呼吸灯,
用按键控制呼吸频率,
单灯或双灯同步等功能.
*/
module RainbowRGB
(input CLK
,input BTN_RST
,output[2:0]RGB
);



endmodule